//Adding anyEdge signal to the transaction class to generate stimulus

class transaction;
  rand bit anyEdge;
  bit risingEdge,fallingEdge;
  
endclass